`default_nettype none

// SDRAM Controller - Winbond W9825G6KH-6 Interface
// 8-state FSM handling initialization, auto-refresh, row activation,
// CAS latency management, and precharge timing for 32 MB synchronous DRAM.
// Supports single-word (32-bit via two 16-bit column accesses) and
// sequential (burst_len>0, pipelined 16-bit column accesses) modes.
// Preserves the internal arbiter interface from sram_controller.sv.
//
// Spec-ref: unit_022_gpu_driver_layer.md `2e395d1315d4c2b1` 2026-02-25

module sdram_controller (
    input  wire         clk,            // 100 MHz system clock (clk_core)
    input  wire         rst_n,          // Active-low synchronous reset

    // ========================================================================
    // Internal memory interface (from arbiter, identical to sram_controller)
    // ========================================================================
    input  wire         req,            // Request signal
    input  wire         we,             // Write enable (1=write, 0=read)
    input  wire [23:0]  addr,           // Byte address (word-aligned, bit 0 unused)
    input  wire [31:0]  wdata,          // Write data (single-word mode)
    output wire [31:0]  rdata,          // Read data (single-word mode, 32-bit assembled)
    output wire         ack,            // Acknowledge (1 cycle pulse)
    output wire         ready,          // Ready for new request

    // Burst interface (from arbiter)
    input  wire [7:0]   burst_len,      // Burst length: 0=single-word, 1-255=sequential (16-bit words)
    input  wire [15:0]  burst_wdata_16, // 16-bit write data for sequential mode
    input  wire         burst_cancel,   // Cancel active burst (from arbiter)
    output wire         burst_data_valid, // Valid 16-bit read data available (sequential read)
    output wire         burst_wdata_req,  // Request next 16-bit write word (sequential write)
    output wire         burst_done,       // Burst transfer complete
    output wire [15:0]  rdata_16,         // 16-bit read data during sequential access

    // ========================================================================
    // External SDRAM interface (directly to W9825G6KH-6 pins)
    // ========================================================================
    // Note: sdram_clk is connected directly from PLL (90-degree phase shifted),
    //       not generated by this module.
    output reg          sdram_cke,      // Clock enable (active high)
    output reg          sdram_csn,      // Chip select (active low)
    output reg          sdram_rasn,     // Row address strobe (active low)
    output reg          sdram_casn,     // Column address strobe (active low)
    output reg          sdram_wen,      // Write enable (active low)
    output reg  [1:0]   sdram_ba,       // Bank address
    output reg  [12:0]  sdram_a,        // Address bus (row: A[12:0], column: A[8:0])
    inout  wire [15:0]  sdram_dq,       // Bidirectional data bus
    output reg  [1:0]   sdram_dqm       // Data mask (upper/lower byte)
);

    // ========================================================================
    // SDRAM Command Encoding
    // {csn, rasn, casn, wen}
    // ========================================================================
    localparam [3:0] CMD_NOP          = 4'b0111;
    localparam [3:0] CMD_ACTIVATE     = 4'b0011;
    localparam [3:0] CMD_READ         = 4'b0101;
    localparam [3:0] CMD_WRITE        = 4'b0100;
    localparam [3:0] CMD_PRECHARGE    = 4'b0010;
    localparam [3:0] CMD_AUTO_REFRESH = 4'b0001;
    localparam [3:0] CMD_LOAD_MODE    = 4'b0000;

    // ========================================================================
    // SDRAM Timing Parameters (100 MHz, W9825G6KH-6)
    // ========================================================================
    localparam INIT_WAIT_CYCLES = 16'd20000;  // 200 us at 100 MHz
    localparam [3:0] T_RCD     = 4'd2;       // RAS to CAS delay (2 cycles)
    localparam [3:0] T_RP      = 4'd2;       // Row precharge time (2 cycles)
    localparam [3:0] T_RC      = 4'd6;       // Row cycle time for auto-refresh (6 cycles)
    localparam [3:0] T_WR      = 4'd2;       // Write recovery time (2 cycles)
    localparam [3:0] T_MRD     = 4'd2;       // Mode register set delay (2 cycles)
    localparam [2:0] CAS_LATENCY = 3'd3;     // CAS latency (3 cycles)
    localparam REFRESH_INTERVAL = 10'd780;    // 781 cycles at 100 MHz (7.81 us per row)

    // Mode register value: CAS latency=3, burst length=1, sequential burst type
    // A[12:10] = reserved (0), A[9] = burst write (0=programmed), A[8:7] = operating mode (00=standard)
    // A[6:4] = CAS latency (011=3), A[3] = burst type (0=sequential), A[2:0] = burst length (000=1)
    localparam [12:0] MODE_REGISTER = 13'b000_0_00_011_0_000;

    // ========================================================================
    // FSM State Definitions (8-state)
    // ========================================================================
    typedef enum logic [2:0] {
        ST_INIT      = 3'd0,
        ST_IDLE      = 3'd1,
        ST_ACTIVATE  = 3'd2,
        ST_READ      = 3'd3,
        ST_WRITE     = 3'd4,
        ST_PRECHARGE = 3'd5,
        ST_REFRESH   = 3'd6,
        ST_DONE      = 3'd7
    } state_t;

    state_t state, next_state;

    // ========================================================================
    // Initialization Sub-State Machine
    // ========================================================================
    typedef enum logic [2:0] {
        INIT_WAIT       = 3'd0,   // 200 us power-up wait
        INIT_PRECHARGE  = 3'd1,   // PRECHARGE ALL
        INIT_PRE_WAIT   = 3'd2,   // Wait tRP
        INIT_REFRESH1   = 3'd3,   // First AUTO REFRESH
        INIT_REFRESH2   = 3'd4,   // Second AUTO REFRESH
        INIT_LOAD_MODE  = 3'd5,   // LOAD MODE REGISTER
        INIT_MODE_WAIT  = 3'd6,   // Wait tMRD
        INIT_COMPLETE   = 3'd7    // Initialization done
    } init_state_t;

    init_state_t init_state;

    // ========================================================================
    // Internal Registers
    // ========================================================================

    // Timing counters
    reg [15:0] init_counter;          // Initialization delay counter
    reg [3:0]  wait_counter;          // General-purpose wait counter for tRCD, tRP, tRC, tWR, tMRD
    reg [9:0]  refresh_timer;         // Auto-refresh interval counter
    reg        refresh_pending;       // Refresh request flag

    // Address decomposition registers
    reg [1:0]  bank_addr;             // Bank address: addr[23:22]
    reg [12:0] row_addr;              // Row address: addr[21:9]
    reg [8:0]  col_addr;              // Column address: addr[8:0] (bit 0 unused for byte alignment)

    // Access control registers
    reg        we_reg;                // Latched write enable
    reg [31:0] wdata_reg;             // Latched write data (single-word mode)
    reg [15:0] rdata_low;             // Low 16 bits of read data (single-word mode)
    reg [31:0] rdata_hold;            // Registered 32-bit read data
    reg [7:0]  burst_count;           // Remaining words in sequential transfer
    reg        burst_mode;            // Sequential transfer active flag
    reg        single_phase;          // 0=low half, 1=high half (single-word mode)

    // Read pipeline tracking for CAS latency
    // For pipelined sequential reads, we issue READ commands every cycle
    // and data arrives CAS_LATENCY cycles later.
    reg [2:0]  read_pipe_count;       // Number of READ commands issued (pipeline fill)
    reg [7:0]  data_remaining;        // Data words still expected from pipeline

    // Write tracking
    reg [7:0]  write_issued;          // Number of WRITE commands issued

    // Data bus control
    reg        dq_oe;                 // Output enable for sdram_dq
    reg [15:0] dq_out;                // Data to drive on sdram_dq

    // Row boundary tracking for sequential access
    reg [8:0]  seq_col;               // Current column for sequential access

    // Precharge-after reason tracking
    reg        precharge_for_refresh; // After precharge, go to REFRESH (else go to DONE)

    // ========================================================================
    // Address alignment check
    // ========================================================================
    // Byte address bit 0 is unused; all SDRAM columns are 16-bit word-aligned.
    // Decomposition uses addr[23:1] only. Declare a wire to suppress the
    // unused-bit warning without a lint pragma.
    wire addr_bit0_unused = addr[0];

    // ========================================================================
    // Bidirectional Data Bus
    // ========================================================================
    assign sdram_dq = dq_oe ? dq_out : 16'bz;
    assign rdata_16 = sdram_dq;

    // ========================================================================
    // SDRAM Command Helper
    // ========================================================================
    // Drives {sdram_csn, sdram_rasn, sdram_casn, sdram_wen} from a 4-bit command
    task automatic set_cmd(input logic [3:0] cmd);
        sdram_csn  = cmd[3];
        sdram_rasn = cmd[2];
        sdram_casn = cmd[1];
        sdram_wen  = cmd[0];
    endtask

    // ========================================================================
    // Output Assignments
    // ========================================================================

    // ready: asserted only in IDLE and not during initialization or refresh
    assign ready = (state == ST_IDLE) && !refresh_pending;

    // ack: single-cycle pulse in DONE state
    assign ack = (state == ST_DONE);

    // burst_done: ack pulse when in burst/sequential mode
    assign burst_done = (state == ST_DONE) && burst_mode;

    // burst_data_valid: valid read data available during sequential read
    // Data is valid when we are in READ state, doing sequential reads,
    // and the CAS latency pipeline has delivered data.
    // Uses read_pipe_count directly (combinational) so that burst_data_valid is asserted on the
    // exact cycle that data first appears on the DQ bus after CAS latency.
    assign burst_data_valid = (state == ST_READ) && burst_mode && !we_reg
                              && (read_pipe_count >= CAS_LATENCY[2:0])
                              && (data_remaining > 8'd0);

    // burst_wdata_req: request next write word during sequential write
    // Asserted after the first WRITE command has been issued (write_issued > 0),
    // indicating the controller has consumed the current word and needs the next.
    // Not asserted on the ACTIVATE->WRITE transition cycle (write_issued still 0)
    // to avoid the arbiter/port advancing data before the first word is captured.
    assign burst_wdata_req = (state == ST_WRITE) && burst_mode && we_reg
                             && (burst_count > 8'd0) && !burst_cancel
                             && (write_issued > 8'd0);

    // rdata: assembled 32-bit word for single-word reads
    // Valid on ack cycle for single-word reads
    assign rdata = rdata_hold;

    // ========================================================================
    // State Machine - Sequential Logic (state register)
    // ========================================================================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= ST_INIT;
        end else begin
            state <= next_state;
        end
    end

    // ========================================================================
    // State Machine - Combinational Logic (next-state)
    // ========================================================================
    always_comb begin
        // Default: stay in current state
        next_state = state;

        case (state)
            ST_INIT: begin
                if (init_state == INIT_COMPLETE) begin
                    next_state = ST_IDLE;
                end
            end

            ST_IDLE: begin
                if (refresh_pending) begin
                    next_state = ST_REFRESH;
                end else if (req) begin
                    next_state = ST_ACTIVATE;
                end
            end

            ST_ACTIVATE: begin
                // Wait tRCD cycles, then go to READ or WRITE
                if (wait_counter == 4'd0) begin
                    if (we_reg) begin
                        next_state = ST_WRITE;
                    end else begin
                        next_state = ST_READ;
                    end
                end
            end

            ST_READ: begin
                // Single-word: wait for both halves to be read
                // Sequential: wait for all pipelined data to arrive
                if (burst_mode) begin
                    // Sequential read: done when all data received or cancelled
                    if (burst_cancel || (data_remaining == 8'd0 && read_pipe_count >= CAS_LATENCY[2:0])) begin
                        next_state = ST_PRECHARGE;
                    end
                end else begin
                    // Single-word read: done when high half data captured
                    // Phase 0: issue READ low, Phase 1: issue READ high
                    // After both READs, wait for CAS latency pipeline to drain
                    if (single_phase && data_remaining == 8'd0 && read_pipe_count >= CAS_LATENCY[2:0]) begin
                        next_state = ST_PRECHARGE;
                    end
                end
            end

            ST_WRITE: begin
                if (burst_mode) begin
                    // Sequential write: done when all writes issued or cancelled
                    if (burst_cancel || burst_count == 8'd0) begin
                        // Need to wait tWR before precharge
                        if (wait_counter == 4'd0) begin
                            next_state = ST_PRECHARGE;
                        end
                    end
                end else begin
                    // Single-word write: done after both halves written + tWR
                    if (single_phase && wait_counter == 4'd0) begin
                        next_state = ST_PRECHARGE;
                    end
                end
            end

            ST_PRECHARGE: begin
                if (wait_counter == 4'd0) begin
                    if (precharge_for_refresh) begin
                        next_state = ST_REFRESH;
                    end else begin
                        next_state = ST_DONE;
                    end
                end
            end

            ST_REFRESH: begin
                if (wait_counter == 4'd0) begin
                    next_state = ST_IDLE;
                end
            end

            ST_DONE: begin
                next_state = ST_IDLE;
            end

            default: begin
                next_state = ST_IDLE;
            end
        endcase
    end

    // ========================================================================
    // Initialization Sub-FSM
    // ========================================================================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            init_state   <= INIT_WAIT;
            init_counter <= INIT_WAIT_CYCLES;
        end else if (state == ST_INIT) begin
            case (init_state)
                INIT_WAIT: begin
                    if (init_counter == 16'd0) begin
                        init_state <= INIT_PRECHARGE;
                    end else begin
                        init_counter <= init_counter - 16'd1;
                    end
                end

                INIT_PRECHARGE: begin
                    // PRECHARGE ALL command issued this cycle (in datapath block)
                    init_state <= INIT_PRE_WAIT;
                end

                INIT_PRE_WAIT: begin
                    // Wait tRP
                    if (wait_counter == 4'd0) begin
                        init_state <= INIT_REFRESH1;
                    end
                end

                INIT_REFRESH1: begin
                    // First AUTO REFRESH issued this cycle
                    // wait_counter loaded with tRC in datapath block
                    if (wait_counter == 4'd0) begin
                        init_state <= INIT_REFRESH2;
                    end
                end

                INIT_REFRESH2: begin
                    // Second AUTO REFRESH issued
                    if (wait_counter == 4'd0) begin
                        init_state <= INIT_LOAD_MODE;
                    end
                end

                INIT_LOAD_MODE: begin
                    // LOAD MODE REGISTER issued this cycle
                    init_state <= INIT_MODE_WAIT;
                end

                INIT_MODE_WAIT: begin
                    // Wait tMRD
                    if (wait_counter == 4'd0) begin
                        init_state <= INIT_COMPLETE;
                    end
                end

                INIT_COMPLETE: begin
                    // Stay here; main FSM transitions to ST_IDLE
                end

                default: begin
                    init_state <= INIT_WAIT;
                end
            endcase
        end
    end

    // ========================================================================
    // Auto-Refresh Timer
    // ========================================================================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            refresh_timer   <= 10'd0;
            refresh_pending <= 1'b0;
        end else begin
            if (state == ST_INIT) begin
                // Don't count during init
                refresh_timer   <= 10'd0;
                refresh_pending <= 1'b0;
            end else if (state == ST_REFRESH && next_state == ST_IDLE) begin
                // Reset timer after refresh completes
                refresh_timer   <= 10'd0;
                refresh_pending <= 1'b0;
            end else begin
                if (refresh_timer >= REFRESH_INTERVAL) begin
                    refresh_pending <= 1'b1;
                end else begin
                    refresh_timer <= refresh_timer + 10'd1;
                end
            end
        end
    end

    // ========================================================================
    // Datapath and SDRAM Signal Control (sequential)
    // ========================================================================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // SDRAM signals: NOP, CKE high, DQM masked
            sdram_cke    <= 1'b1;
            sdram_csn    <= 1'b1;
            sdram_rasn   <= 1'b1;
            sdram_casn   <= 1'b1;
            sdram_wen    <= 1'b1;
            sdram_ba     <= 2'b00;
            sdram_a      <= 13'b0;
            sdram_dqm    <= 2'b11;    // Masked during reset
            dq_oe        <= 1'b0;
            dq_out       <= 16'b0;

            // Internal registers
            we_reg            <= 1'b0;
            wdata_reg         <= 32'b0;
            rdata_low         <= 16'b0;
            rdata_hold        <= 32'b0;
            burst_count       <= 8'b0;
            burst_mode        <= 1'b0;
            single_phase      <= 1'b0;
            wait_counter      <= 4'b0;
            read_pipe_count   <= 3'b0;
            data_remaining    <= 8'b0;
            write_issued      <= 8'b0;
            bank_addr         <= 2'b0;
            row_addr          <= 13'b0;
            col_addr          <= 9'b0;
            seq_col           <= 9'b0;
            precharge_for_refresh <= 1'b0;

        end else begin

            case (state)
                // ============================================================
                // INIT: Power-up initialization sequence
                // ============================================================
                ST_INIT: begin
                    sdram_cke <= 1'b1;
                    sdram_dqm <= 2'b11;  // Masked during init
                    dq_oe     <= 1'b0;

                    case (init_state)
                        INIT_WAIT: begin
                            // NOP during power-up wait
                            set_cmd(CMD_NOP);
                        end

                        INIT_PRECHARGE: begin
                            // PRECHARGE ALL (A10=1)
                            set_cmd(CMD_PRECHARGE);
                            sdram_a    <= 13'b0_0100_0000_0000; // A10=1 for all banks
                            sdram_ba   <= 2'b00;
                            wait_counter <= T_RP - 4'd1;
                        end

                        INIT_PRE_WAIT: begin
                            set_cmd(CMD_NOP);
                            if (wait_counter > 4'd0) begin
                                wait_counter <= wait_counter - 4'd1;
                            end
                        end

                        INIT_REFRESH1: begin
                            if (wait_counter == T_RC - 4'd1) begin
                                // Issue AUTO REFRESH on entry
                                set_cmd(CMD_AUTO_REFRESH);
                            end else begin
                                set_cmd(CMD_NOP);
                            end
                            if (wait_counter > 4'd0) begin
                                wait_counter <= wait_counter - 4'd1;
                            end else begin
                                // Reload counter for second refresh
                                wait_counter <= T_RC - 4'd1;
                            end
                        end

                        INIT_REFRESH2: begin
                            if (wait_counter == T_RC - 4'd1) begin
                                // Issue second AUTO REFRESH on entry
                                set_cmd(CMD_AUTO_REFRESH);
                            end else begin
                                set_cmd(CMD_NOP);
                            end
                            if (wait_counter > 4'd0) begin
                                wait_counter <= wait_counter - 4'd1;
                            end
                        end

                        INIT_LOAD_MODE: begin
                            // LOAD MODE REGISTER
                            set_cmd(CMD_LOAD_MODE);
                            sdram_a  <= MODE_REGISTER;
                            sdram_ba <= 2'b00;
                            wait_counter <= T_MRD - 4'd1;
                        end

                        INIT_MODE_WAIT: begin
                            set_cmd(CMD_NOP);
                            if (wait_counter > 4'd0) begin
                                wait_counter <= wait_counter - 4'd1;
                            end
                        end

                        INIT_COMPLETE: begin
                            set_cmd(CMD_NOP);
                            sdram_dqm <= 2'b00;  // Unmask for normal operation
                        end

                        default: begin
                            set_cmd(CMD_NOP);
                        end
                    endcase
                end

                // ============================================================
                // IDLE: Ready for requests; check refresh
                // ============================================================
                ST_IDLE: begin
                    set_cmd(CMD_NOP);
                    dq_oe     <= 1'b0;
                    sdram_dqm <= 2'b00;
                    precharge_for_refresh <= 1'b0;

                    if (refresh_pending && !req) begin
                        // Refresh will be handled in next state
                    end else if (req) begin
                        // Latch request parameters
                        we_reg     <= we;
                        wdata_reg  <= wdata;
                        burst_mode <= (burst_len > 8'd0);
                        burst_count <= burst_len;
                        single_phase <= 1'b0;
                        read_pipe_count   <= 3'b0;
                        data_remaining    <= 8'b0;
                        write_issued      <= 8'b0;

                        // Address decomposition:
                        // addr[23:0] is a byte address into 32 MB space
                        // Bit 0 is unused (word-aligned)
                        // For SDRAM: bank = addr[23:22], row = addr[21:9], col = addr[8:1]
                        // But our column width is 9 bits (512 columns), so:
                        // bank = addr[23:22]
                        // row  = addr[21:9]
                        // col  = addr[8:1] with bit 0 of column always 0 for 16-bit access
                        bank_addr <= addr[23:22];
                        row_addr  <= addr[21:9];
                        col_addr  <= {addr[8:1], 1'b0}; // Column address (9 bits, aligned)
                        seq_col   <= {addr[8:1], 1'b0};
                    end
                end

                // ============================================================
                // ACTIVATE: Open row in target bank
                // ============================================================
                ST_ACTIVATE: begin
                    if (wait_counter == T_RCD) begin
                        // First cycle: issue ACTIVATE command
                        set_cmd(CMD_ACTIVATE);
                        sdram_ba <= bank_addr;
                        sdram_a  <= row_addr;
                        wait_counter <= wait_counter - 4'd1;
                    end else if (wait_counter > 4'd0) begin
                        // Waiting tRCD
                        set_cmd(CMD_NOP);
                        wait_counter <= wait_counter - 4'd1;
                    end else begin
                        // tRCD elapsed, transition to READ or WRITE
                        set_cmd(CMD_NOP);
                    end
                end

                // ============================================================
                // READ: Issue READ commands and capture data after CAS latency
                // ============================================================
                ST_READ: begin
                    if (burst_mode) begin
                        // ----- Sequential Read -----
                        // Issue pipelined READ commands to consecutive columns
                        // Data arrives CAS_LATENCY cycles after each READ

                        // Determine if we are issuing a READ and/or receiving data
                        // this cycle, then compute a single data_remaining update
                        // to avoid conflicting NBA assignments.

                        if (burst_count > 8'd0 && !burst_cancel) begin
                            // Issue next READ command
                            set_cmd(CMD_READ);
                            sdram_ba <= bank_addr;
                            sdram_a  <= {4'b0, seq_col}; // A10=0 (no auto-precharge)
                            seq_col  <= seq_col + 9'd1;
                            burst_count <= burst_count - 8'd1;
                            read_pipe_count <= (read_pipe_count < CAS_LATENCY[2:0]) ?
                                               read_pipe_count + 3'd1 : read_pipe_count;

                            // data_remaining: +1 for issued READ, -1 if data also arriving
                            if (read_pipe_count >= CAS_LATENCY[2:0] && data_remaining > 8'd0) begin
                                // Both issuing and receiving: net change is 0
                                // data_remaining stays the same (no assignment needed)
                            end else begin
                                data_remaining <= data_remaining + 8'd1;
                            end
                        end else begin
                            // No more READs to issue; wait for pipeline to drain
                            set_cmd(CMD_NOP);
                            if (read_pipe_count < CAS_LATENCY[2:0]) begin
                                read_pipe_count <= read_pipe_count + 3'd1;
                            end

                            // Data arrives CAS_LATENCY cycles after first READ
                            if (read_pipe_count >= CAS_LATENCY[2:0] && data_remaining > 8'd0) begin
                                data_remaining <= data_remaining - 8'd1;
                            end
                        end

                        dq_oe <= 1'b0;

                    end else begin
                        // ----- Single-Word Read -----
                        // Two sequential READ commands: low half then high half
                        if (!single_phase) begin
                            if (read_pipe_count == 3'd0) begin
                                // Issue READ for low half
                                set_cmd(CMD_READ);
                                sdram_ba <= bank_addr;
                                sdram_a  <= {4'b0, col_addr}; // A10=0
                                read_pipe_count <= 3'd1;
                                data_remaining  <= 8'd1;
                            end else if (read_pipe_count < CAS_LATENCY[2:0]) begin
                                set_cmd(CMD_NOP);
                                read_pipe_count <= read_pipe_count + 3'd1;
                            end else begin
                                // CAS latency elapsed; latch low data
                                set_cmd(CMD_NOP);
                                rdata_low <= sdram_dq;
                                data_remaining  <= 8'd0;
                                // Move to high half
                                single_phase    <= 1'b1;
                                read_pipe_count <= 3'd0;
                            end
                        end else begin
                            if (read_pipe_count == 3'd0) begin
                                // Issue READ for high half (col + 1)
                                set_cmd(CMD_READ);
                                sdram_ba <= bank_addr;
                                sdram_a  <= {4'b0, col_addr + 9'd1}; // A10=0
                                read_pipe_count <= 3'd1;
                                data_remaining  <= 8'd1;
                            end else if (read_pipe_count < CAS_LATENCY[2:0]) begin
                                set_cmd(CMD_NOP);
                                read_pipe_count <= read_pipe_count + 3'd1;
                            end else begin
                                // CAS latency elapsed; latch high data and assemble
                                set_cmd(CMD_NOP);
                                rdata_hold <= {sdram_dq, rdata_low};
                                data_remaining <= 8'd0;
                            end
                        end

                        dq_oe <= 1'b0;
                    end
                end

                // ============================================================
                // WRITE: Issue WRITE commands with data
                // ============================================================
                ST_WRITE: begin
                    if (burst_mode) begin
                        // ----- Sequential Write -----
                        if (burst_count > 8'd0 && !burst_cancel) begin
                            // Issue WRITE command with data
                            set_cmd(CMD_WRITE);
                            sdram_ba <= bank_addr;
                            sdram_a  <= {4'b0, seq_col}; // A10=0
                            dq_oe    <= 1'b1;
                            dq_out   <= burst_wdata_16;
                            seq_col  <= seq_col + 9'd1;
                            burst_count  <= burst_count - 8'd1;
                            write_issued <= write_issued + 8'd1;
                            wait_counter <= T_WR; // Reset tWR counter after each write
                        end else begin
                            // All writes issued or cancelled; wait tWR
                            set_cmd(CMD_NOP);
                            dq_oe <= 1'b0;
                            if (wait_counter > 4'd0) begin
                                wait_counter <= wait_counter - 4'd1;
                            end
                        end

                    end else begin
                        // ----- Single-Word Write -----
                        if (!single_phase) begin
                            // Write low half
                            set_cmd(CMD_WRITE);
                            sdram_ba <= bank_addr;
                            sdram_a  <= {4'b0, col_addr}; // A10=0
                            dq_oe    <= 1'b1;
                            dq_out   <= wdata_reg[15:0];
                            single_phase <= 1'b1;
                            wait_counter <= T_WR; // Will be refreshed after high write
                        end else begin
                            if (write_issued == 8'd0) begin
                                // Write high half (col + 1)
                                set_cmd(CMD_WRITE);
                                sdram_ba <= bank_addr;
                                sdram_a  <= {4'b0, col_addr + 9'd1}; // A10=0
                                dq_oe    <= 1'b1;
                                dq_out   <= wdata_reg[31:16];
                                write_issued <= 8'd1;
                                wait_counter <= T_WR; // Start tWR after last write
                            end else begin
                                // Wait tWR
                                set_cmd(CMD_NOP);
                                dq_oe <= 1'b0;
                                if (wait_counter > 4'd0) begin
                                    wait_counter <= wait_counter - 4'd1;
                                end
                            end
                        end
                    end
                end

                // ============================================================
                // PRECHARGE: Close active row
                // ============================================================
                ST_PRECHARGE: begin
                    if (wait_counter == T_RP) begin
                        // First cycle: issue PRECHARGE command
                        set_cmd(CMD_PRECHARGE);
                        sdram_ba <= bank_addr;
                        sdram_a  <= precharge_for_refresh ? 13'b0_0100_0000_0000 : 13'b0; // A10=1 for all-bank if refresh
                        dq_oe    <= 1'b0;
                        wait_counter <= wait_counter - 4'd1;
                    end else if (wait_counter > 4'd0) begin
                        set_cmd(CMD_NOP);
                        wait_counter <= wait_counter - 4'd1;
                    end else begin
                        set_cmd(CMD_NOP);
                    end
                end

                // ============================================================
                // REFRESH: Execute AUTO REFRESH
                // ============================================================
                ST_REFRESH: begin
                    if (wait_counter == T_RC - 4'd1) begin
                        // First cycle: issue AUTO REFRESH
                        set_cmd(CMD_AUTO_REFRESH);
                        wait_counter <= wait_counter - 4'd1;
                    end else if (wait_counter > 4'd0) begin
                        set_cmd(CMD_NOP);
                        wait_counter <= wait_counter - 4'd1;
                    end else begin
                        set_cmd(CMD_NOP);
                    end
                end

                // ============================================================
                // DONE: Acknowledge completion
                // ============================================================
                ST_DONE: begin
                    set_cmd(CMD_NOP);
                    dq_oe     <= 1'b0;
                    burst_mode <= 1'b0;
                end

                default: begin
                    set_cmd(CMD_NOP);
                    dq_oe <= 1'b0;
                end
            endcase

            // ================================================================
            // Wait counter initialization on state transitions
            // ================================================================
            // Load wait counter when transitioning to states that need it
            if (state != next_state) begin
                case (next_state)
                    ST_ACTIVATE: begin
                        wait_counter <= T_RCD;
                    end
                    ST_PRECHARGE: begin
                        wait_counter <= T_RP;
                        // Determine where to go after precharge
                        precharge_for_refresh <= refresh_pending;
                    end
                    ST_REFRESH: begin
                        wait_counter <= T_RC - 4'd1;
                    end
                    default: begin
                        // No explicit wait counter load needed
                    end
                endcase
            end
        end
    end

endmodule
