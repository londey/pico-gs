// Testbench for Triangle Rasterizer (Incremental Interpolation, DD-024)
// Tests basic triangle rasterization with edge functions, fragment output bus,
// derivative precomputation, and incremental attribute interpolation.
// Includes parametric bounding-box clamping tests for multiple surface sizes.
//
// Verification reference: VER-001 (Rasterizer Unit Testbench)
// Spec-ref: unit_005_rasterizer.md `0000000000000000` 1970-01-01

`timescale 1ns/1ps

module tb_rasterizer;
    import fp_types_pkg::*;

    // Clock and reset
    reg clk;
    reg rst_n;

    // Triangle input
    reg         tri_valid;
    wire        tri_ready;

    reg [15:0]  v0_x, v0_y, v0_z;
    reg [31:0]  v0_color0, v0_color1;
    reg [31:0]  v0_uv0, v0_uv1;
    reg [15:0]  v0_q;

    reg [15:0]  v1_x, v1_y, v1_z;
    reg [31:0]  v1_color0, v1_color1;
    reg [31:0]  v1_uv0, v1_uv1;
    reg [15:0]  v1_q;

    reg [15:0]  v2_x, v2_y, v2_z;
    reg [31:0]  v2_color0, v2_color1;
    reg [31:0]  v2_uv0, v2_uv1;
    reg [15:0]  v2_q;

    // Inverse area
    reg [15:0]  inv_area;

    // Fragment output bus
    wire        frag_valid;
    reg         frag_ready;
    wire [9:0]  frag_x;
    wire [9:0]  frag_y;
    wire [15:0] frag_z;
    wire [63:0] frag_color0;
    wire [63:0] frag_color1;
    wire [31:0] frag_uv0;
    wire [31:0] frag_uv1;
    wire [15:0] frag_q;

    // Framebuffer surface dimensions (from FB_CONFIG register)
    reg [3:0]   fb_width_log2;
    reg [3:0]   fb_height_log2;

    // Test result tracking
    integer test_pass_count = 0;
    integer test_fail_count = 0;

    // Instantiate DUT
    rasterizer dut (
        .clk(clk),
        .rst_n(rst_n),
        .tri_valid(tri_valid),
        .tri_ready(tri_ready),

        .v0_x(v0_x), .v0_y(v0_y), .v0_z(v0_z),
        .v0_color0(v0_color0), .v0_color1(v0_color1),
        .v0_uv0(v0_uv0), .v0_uv1(v0_uv1), .v0_q(v0_q),

        .v1_x(v1_x), .v1_y(v1_y), .v1_z(v1_z),
        .v1_color0(v1_color0), .v1_color1(v1_color1),
        .v1_uv0(v1_uv0), .v1_uv1(v1_uv1), .v1_q(v1_q),

        .v2_x(v2_x), .v2_y(v2_y), .v2_z(v2_z),
        .v2_color0(v2_color0), .v2_color1(v2_color1),
        .v2_uv0(v2_uv0), .v2_uv1(v2_uv1), .v2_q(v2_q),

        .inv_area(inv_area),

        .frag_valid(frag_valid),
        .frag_ready(frag_ready),
        .frag_x(frag_x),
        .frag_y(frag_y),
        .frag_z(frag_z),
        .frag_color0(frag_color0),
        .frag_color1(frag_color1),
        .frag_uv0(frag_uv0),
        .frag_uv1(frag_uv1),
        .frag_q(frag_q),

        .fb_width_log2(fb_width_log2),
        .fb_height_log2(fb_height_log2)
    );

    // Clock generation (100 MHz system clock)
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // ========================================================================
    // Helper task: submit a triangle and wait for rasterization to complete
    // ========================================================================
    task submit_triangle_and_wait;
        begin
            tri_valid = 1;
            @(posedge clk);
            wait(tri_ready == 0);  // Wait for rasterizer to accept
            tri_valid = 0;
            // Wait for rasterization to complete
            wait(tri_ready == 1);
        end
    endtask

    // ========================================================================
    // Helper task: check parametric bounding-box clamping
    // ========================================================================
    task check_bbox_clamp(
        input [3:0] width_log2,
        input [3:0] height_log2,
        input string test_label
    );
        reg [9:0] max_x_bound;
        reg [9:0] max_y_bound;
        begin
            max_x_bound = (10'd1 << width_log2) - 10'd1;
            max_y_bound = (10'd1 << height_log2) - 10'd1;

            if (dut.bbox_max_x <= max_x_bound) begin
                $display("  PASS: %s bbox_max_x=%0d <= %0d", test_label, dut.bbox_max_x, max_x_bound);
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("  FAIL: %s bbox_max_x=%0d > %0d", test_label, dut.bbox_max_x, max_x_bound);
                test_fail_count = test_fail_count + 1;
            end

            if (dut.bbox_max_y <= max_y_bound) begin
                $display("  PASS: %s bbox_max_y=%0d <= %0d", test_label, dut.bbox_max_y, max_y_bound);
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("  FAIL: %s bbox_max_y=%0d > %0d", test_label, dut.bbox_max_y, max_y_bound);
                test_fail_count = test_fail_count + 1;
            end
        end
    endtask

    // ========================================================================
    // Helper task: set default vertex attributes (zero UV, color1, Q)
    // ========================================================================
    task set_default_attrs;
        begin
            v0_color1 = 32'h00000000;
            v0_uv0 = 32'h00000000;
            v0_uv1 = 32'h00000000;
            v0_q = 16'h1000;  // Q = 1.0 in Q3.12

            v1_color1 = 32'h00000000;
            v1_uv0 = 32'h00000000;
            v1_uv1 = 32'h00000000;
            v1_q = 16'h1000;

            v2_color1 = 32'h00000000;
            v2_uv0 = 32'h00000000;
            v2_uv1 = 32'h00000000;
            v2_q = 16'h1000;
        end
    endtask

    // ========================================================================
    // Fragment counter and monitor
    // ========================================================================
    integer pixel_count = 0;
    integer total_frag_count = 0;

    always @(posedge clk) begin
        if (frag_valid && frag_ready) begin
            pixel_count = pixel_count + 1;
            total_frag_count = total_frag_count + 1;

            // Debug first few pixels per triangle
            if (pixel_count <= 3) begin
                $display("  Fragment %0d: x=%0d y=%0d z=0x%04x color0=0x%016x",
                         pixel_count, frag_x, frag_y, frag_z, frag_color0);
            end
        end
    end

    // ========================================================================
    // Interpolation reference model (incremental stepping, DD-024)
    // ========================================================================
    // Replicates the rasterizer's derivative precomputation and output
    // promotion logic in the testbench for comparison.  Uses the same
    // fixed-point widths and truncation rules as the RTL.

    // Compute a single 8-bit-channel derivative (dx or dy) using the same
    // formula as the rasterizer: raw = d10*coeff_A1 + d20*coeff_A2,
    // then scaled = (raw * inv_area_val) >>> 16.
    function automatic signed [31:0] ref_deriv_8bit(
        input [7:0] f0, input [7:0] f1, input [7:0] f2,
        input signed [10:0] coeff1, input signed [10:0] coeff2,
        input [15:0] inv_area_val
    );
        reg signed [8:0]  d10, d20;
        reg signed [20:0] raw;
        reg signed [36:0] scl;
        begin
            d10 = $signed({1'b0, f1}) - $signed({1'b0, f0});
            d20 = $signed({1'b0, f2}) - $signed({1'b0, f0});
            raw = (d10 * coeff1) + (d20 * coeff2);
            scl = raw * $signed({1'b0, inv_area_val});
            ref_deriv_8bit = scl >>> 16;
        end
    endfunction

    // Compute a single 16-bit-channel derivative (dx or dy) for Z (unsigned
    // origin), UV (signed), or Q (unsigned origin).
    function automatic signed [31:0] ref_deriv_16bit(
        input signed [16:0] d10, input signed [16:0] d20,
        input signed [10:0] coeff1, input signed [10:0] coeff2,
        input [15:0] inv_area_val
    );
        reg signed [28:0] raw;
        reg signed [44:0] scl;
        begin
            raw = (d10 * coeff1) + (d20 * coeff2);
            scl = raw * $signed({1'b0, inv_area_val});
            ref_deriv_16bit = scl >>> 16;
        end
    endfunction

    // Promote an 8.16 accumulator to Q4.12, matching the RTL clamp logic.
    function automatic [15:0] ref_promote_8bit(input signed [31:0] acc);
        begin
            if (acc[31]) begin
                ref_promote_8bit = 16'h0000;
            end else if (acc[31:24] != 8'd0) begin
                ref_promote_8bit = {4'b0, 8'hFF, 4'hF};
            end else begin
                ref_promote_8bit = {4'b0, acc[23:16], acc[23:20]};
            end
        end
    endfunction

    // Promote Z accumulator to 16-bit output, matching the RTL clamp logic.
    function automatic [15:0] ref_promote_z(input signed [31:0] acc);
        begin
            if (acc[31]) begin
                ref_promote_z = 16'h0000;
            end else begin
                ref_promote_z = acc[31:16];
            end
        end
    endfunction

    // ========================================================================
    // Test sequence
    // ========================================================================
    initial begin
        $dumpfile("rasterizer.vcd");
        $dumpvars(0, tb_rasterizer);

        // Initialize
        rst_n = 0;
        tri_valid = 0;
        frag_ready = 1;  // Always accept fragments by default

        // Default surface dimensions: 512x512 (VER-001 precondition)
        fb_width_log2  = 4'd9;
        fb_height_log2 = 4'd9;

        // Default attributes
        set_default_attrs;

        #100;
        rst_n = 1;
        #100;

        $display("=== Testing Triangle Rasterizer (Incremental Interpolation) ===\n");

        // ====================================================================
        // Test 1: Small triangle at origin (512x512 surface)
        // Verifies: edge function coefficients, fragment emission, bbox
        // (VER-001 steps 1 and 3)
        // ====================================================================
        $display("Test 1: Small triangle (10,10) -> (50,10) -> (30,40) [512x512 surface]");
        fb_width_log2  = 4'd9;
        fb_height_log2 = 4'd9;
        pixel_count = 0;

        // Vertex 0: (10, 10) in 12.4 fixed point = 10 << 4 = 160
        v0_x = 16'd160;
        v0_y = 16'd160;
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;  // Red (RGBA8888)
        set_default_attrs;

        // Vertex 1: (50, 10)
        v1_x = 16'd800;  // 50 << 4
        v1_y = 16'd160;
        v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;  // Green

        // Vertex 2: (30, 40)
        v2_x = 16'd480;  // 30 << 4
        v2_y = 16'd640;  // 40 << 4
        v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;  // Blue

        // inv_area = 65536/1200 ~ 55 = 0x0037
        inv_area = 16'h0037;

        submit_triangle_and_wait;
        $display("  Triangle rasterization completed at time %0t, fragments=%0d", $time, pixel_count);

        // Check that bbox is within 512x512 bounds
        check_bbox_clamp(4'd9, 4'd9, "Test1-within-bounds");

        // Verify fragments were emitted
        if (pixel_count > 0) begin
            $display("  PASS: Fragment count > 0 (%0d fragments)", pixel_count);
            test_pass_count = test_pass_count + 1;
        end else begin
            $display("  FAIL: No fragments emitted");
            test_fail_count = test_fail_count + 1;
        end

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 2a: Bounding-box clamping on 512x512 surface (VER-001 step 2a)
        // ====================================================================
        $display("\nTest 2a: Bbox clamping on 512x512 surface -- triangle out of bounds");
        fb_width_log2  = 4'd9;
        fb_height_log2 = 4'd9;
        pixel_count = 0;

        v0_x = 16'd8080;  // 505 << 4
        v0_y = 16'd8080;
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;
        set_default_attrs;

        v1_x = 16'd8320;  // 520 << 4
        v1_y = 16'd8080;
        v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;

        v2_x = 16'd8160;  // 510 << 4
        v2_y = 16'd8320;  // 520 << 4
        v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;

        inv_area = 16'h0200;

        submit_triangle_and_wait;
        $display("  Triangle rasterization completed at time %0t", $time);
        check_bbox_clamp(4'd9, 4'd9, "Test2a-512x512-clamped");

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 2a-within: Fully within 512x512 bounds
        // ====================================================================
        $display("\nTest 2a-within: Triangle fully within 512x512 bounds");
        fb_width_log2  = 4'd9;
        fb_height_log2 = 4'd9;
        pixel_count = 0;

        v0_x = 16'd1600;  // 100 << 4
        v0_y = 16'd1600;
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;
        set_default_attrs;

        v1_x = 16'd1920;  // 120 << 4
        v1_y = 16'd1600;
        v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;

        v2_x = 16'd1760;  // 110 << 4
        v2_y = 16'd1920;  // 120 << 4
        v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;

        inv_area = 16'h0200;

        submit_triangle_and_wait;
        $display("  Triangle rasterization completed at time %0t", $time);
        check_bbox_clamp(4'd9, 4'd9, "Test2a-within-512x512");

        // Verify bbox matches raw vertex extents (not clamped)
        if (dut.bbox_min_x == 10'd100 && dut.bbox_max_x == 10'd120 &&
            dut.bbox_min_y == 10'd100 && dut.bbox_max_y == 10'd120) begin
            $display("  PASS: bbox matches raw vertex extents [100,120] x [100,120]");
            test_pass_count = test_pass_count + 1;
        end else begin
            $display("  FAIL: bbox does not match expected raw extents");
            $display("        got [%0d,%0d] x [%0d,%0d], expected [100,120] x [100,120]",
                     dut.bbox_min_x, dut.bbox_max_x, dut.bbox_min_y, dut.bbox_max_y);
            test_fail_count = test_fail_count + 1;
        end

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 2b: Bounding-box clamping on 256x256 surface (VER-001 step 2b)
        // ====================================================================
        $display("\nTest 2b: Bbox clamping on 256x256 surface -- triangle out of bounds");
        fb_width_log2  = 4'd8;
        fb_height_log2 = 4'd8;
        pixel_count = 0;

        v0_x = 16'd4000;  // 250 << 4
        v0_y = 16'd4000;
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;
        set_default_attrs;

        v1_x = 16'd4320;  // 270 << 4
        v1_y = 16'd4000;
        v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;

        v2_x = 16'd4160;  // 260 << 4
        v2_y = 16'd4320;  // 270 << 4
        v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;

        inv_area = 16'h0200;

        submit_triangle_and_wait;
        $display("  Triangle rasterization completed at time %0t", $time);
        check_bbox_clamp(4'd8, 4'd8, "Test2b-256x256-clamped");

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 2b-within: Fully within 256x256 bounds
        // ====================================================================
        $display("\nTest 2b-within: Triangle fully within 256x256 bounds");
        fb_width_log2  = 4'd8;
        fb_height_log2 = 4'd8;
        pixel_count = 0;

        v0_x = 16'd800;   // 50 << 4
        v0_y = 16'd800;
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;
        set_default_attrs;

        v1_x = 16'd1120;  // 70 << 4
        v1_y = 16'd800;
        v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;

        v2_x = 16'd960;   // 60 << 4
        v2_y = 16'd1120;  // 70 << 4
        v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;

        inv_area = 16'h0200;

        submit_triangle_and_wait;
        $display("  Triangle rasterization completed at time %0t", $time);
        check_bbox_clamp(4'd8, 4'd8, "Test2b-within-256x256");

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 3: Degenerate triangle -- zero-area collinear vertices
        // (VER-001 step 6)
        // ====================================================================
        $display("\nTest 3: Degenerate triangle -- collinear vertices [512x512 surface]");
        fb_width_log2  = 4'd9;
        fb_height_log2 = 4'd9;
        pixel_count = 0;

        v0_x = 16'd800;   // 50 << 4
        v0_y = 16'd1600;  // 100 << 4
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;
        set_default_attrs;

        v1_x = 16'd1600;  // 100 << 4
        v1_y = 16'd1600;
        v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;

        v2_x = 16'd2400;  // 150 << 4
        v2_y = 16'd1600;
        v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;

        inv_area = 16'h0000;

        submit_triangle_and_wait;
        $display("  Degenerate triangle completed at time %0t, fragments=%0d", $time, pixel_count);

        check_bbox_clamp(4'd9, 4'd9, "Test3-degenerate");

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 3b: Degenerate triangle -- fully off-screen (VER-001 step 6)
        // All vertices outside the configured surface bounds; bounding box
        // clamp should result in an empty region, emitting zero fragments.
        // ====================================================================
        $display("\nTest 3b: Degenerate triangle -- fully off-screen [256x256 surface]");
        fb_width_log2  = 4'd8;
        fb_height_log2 = 4'd8;
        pixel_count = 0;

        // All three vertices at pixel coordinates well above 255
        v0_x = 16'd8160;  // 510 << 4
        v0_y = 16'd8160;
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;
        set_default_attrs;

        v1_x = 16'd8320;  // 520 << 4
        v1_y = 16'd8160;
        v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;

        v2_x = 16'd8240;  // 515 << 4
        v2_y = 16'd8320;  // 520 << 4
        v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;

        inv_area = 16'h0200;

        submit_triangle_and_wait;
        $display("  Off-screen triangle completed at time %0t, fragments=%0d", $time, pixel_count);

        // Verify bounding box was clamped to surface bounds
        check_bbox_clamp(4'd8, 4'd8, "Test3b-offscreen-256x256");

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 4: Fragment output bus back-pressure (VER-001 step 5)
        // After starting a triangle render, assert frag_ready=0 for 5 cycles
        // while fragments are being generated.  Verify no frag_valid
        // transitions during stall, then resume and count total fragments.
        // ====================================================================
        $display("\nTest 4: Fragment output bus back-pressure test");
        fb_width_log2  = 4'd9;
        fb_height_log2 = 4'd9;
        pixel_count = 0;

        // Small triangle that definitely has inside pixels
        v0_x = 16'd320;   // 20 << 4
        v0_y = 16'd320;
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;
        set_default_attrs;

        v1_x = 16'd640;   // 40 << 4
        v1_y = 16'd320;
        v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;

        v2_x = 16'd480;   // 30 << 4
        v2_y = 16'd640;   // 40 << 4
        v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;

        inv_area = 16'h0200;

        // Deassert ready to test back-pressure
        frag_ready = 0;

        tri_valid = 1;
        @(posedge clk);
        wait(tri_ready == 0);
        tri_valid = 0;

        // Wait for rasterizer to reach INTERPOLATE (DD-025 handshake).
        // Need enough cycles for setup (SETUP -> SETUP_2 -> SETUP_3 ->
        // ITER_START -> INIT_E1 -> INIT_E2 -> EDGE_TEST -> INTERPOLATE).
        repeat(20) @(posedge clk);

        // If frag_valid is asserted and we haven't accepted, pixel_count should be 0
        if (pixel_count == 0 && frag_valid) begin
            $display("  PASS: Back-pressure held -- frag_valid=1 but no fragments consumed");
            test_pass_count = test_pass_count + 1;
        end else if (pixel_count == 0) begin
            // Triangle might not have inside pixels at this point, or setup not done
            $display("  INFO: frag_valid=%0d, pixel_count=%0d (may need more cycles)", frag_valid, pixel_count);
        end else begin
            $display("  FAIL: Fragments consumed while frag_ready=0 (pixel_count=%0d)", pixel_count);
            test_fail_count = test_fail_count + 1;
        end

        // Hold back-pressure for 5 more cycles and verify no frag_valid transitions
        begin : bp_stall_check
            integer bp_cycle;
            reg frag_valid_snapshot;
            integer bp_fail;
            frag_valid_snapshot = frag_valid;
            bp_fail = 0;
            for (bp_cycle = 0; bp_cycle < 5; bp_cycle = bp_cycle + 1) begin
                @(posedge clk);
                // During back-pressure, frag_valid should stay high (stalled) and
                // pixel_count should not increase
                if (pixel_count != 0) begin
                    bp_fail = 1;
                end
            end
            if (bp_fail == 0) begin
                $display("  PASS: No fragments consumed during 5-cycle back-pressure stall");
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("  FAIL: Fragments consumed during back-pressure stall");
                test_fail_count = test_fail_count + 1;
            end
        end

        // Record pre-resume count
        begin : bp_resume
            integer pre_resume_count;
            pre_resume_count = pixel_count;

            // Re-assert ready and let rasterization complete
            frag_ready = 1;
            wait(tri_ready == 1);
            $display("  Back-pressure test completed, total fragments=%0d", pixel_count);

            if (pixel_count > pre_resume_count) begin
                $display("  PASS: Fragments emitted after ready re-asserted (%0d fragments)", pixel_count);
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("  FAIL: No fragments emitted after ready re-asserted");
                test_fail_count = test_fail_count + 1;
            end
        end

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 5: Q4.12 UV interpolation with wrapping range (VER-001 step 7)
        // Verifies UV values > 1.0 and negative UV are handled correctly.
        // Q4.12: 1.0 = 0x1000, 2.0 = 0x2000, -1.0 = 0xF000
        // ====================================================================
        $display("\nTest 5: Q4.12 UV interpolation -- wrapping range");
        fb_width_log2  = 4'd9;
        fb_height_log2 = 4'd9;
        pixel_count = 0;

        // Small triangle: (10,10) -> (20,10) -> (15,20)
        v0_x = 16'd160;   // 10 << 4
        v0_y = 16'd160;
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;
        v0_color1 = 32'h00000000;
        // UV0: U=0.0, V=0.0 in Q4.12
        v0_uv0 = {16'h0000, 16'h0000};
        v0_uv1 = 32'h00000000;
        v0_q = 16'h1000;

        v1_x = 16'd320;   // 20 << 4
        v1_y = 16'd160;
        v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;
        v1_color1 = 32'h00000000;
        // UV0: U=2.0, V=0.0 -- wraps past 1.0
        v1_uv0 = {16'h2000, 16'h0000};
        v1_uv1 = 32'h00000000;
        v1_q = 16'h1000;

        v2_x = 16'd240;   // 15 << 4
        v2_y = 16'd320;   // 20 << 4
        v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;
        v2_color1 = 32'h00000000;
        // UV0: U=-1.0, V=2.0 -- negative U, wrapping V
        v2_uv0 = {16'hF000, 16'h2000};
        v2_uv1 = 32'h00000000;
        v2_q = 16'h1000;

        inv_area = 16'h0200;

        submit_triangle_and_wait;
        $display("  Q4.12 UV test completed at time %0t, fragments=%0d", $time, pixel_count);

        if (pixel_count > 0) begin
            $display("  PASS: Fragments emitted with Q4.12 UV wrapping range (%0d fragments)", pixel_count);
            test_pass_count = test_pass_count + 1;
        end else begin
            $display("  FAIL: No fragments emitted");
            test_fail_count = test_fail_count + 1;
        end

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 6: Verify no SDRAM ports exist (VER-001 verification criterion 3)
        // ====================================================================
        $display("\nTest 6: Verify fragment output bus interface (no SDRAM ports)");
        // This is a structural check -- the fact that the DUT compiles with
        // frag_valid/frag_ready and without fb_req/zb_req proves the interface.
        $display("  PASS: DUT compiled with fragment output bus (no SDRAM ports)");
        test_pass_count = test_pass_count + 1;

        // ====================================================================
        // Test 7: Incremental interpolation accuracy (VER-001 step 4)
        // Uses a known triangle with distinct color, Z, UV, and Q values.
        // Computes reference derivatives and initial values using the same
        // formula as the rasterizer, then checks the first emitted fragment
        // for a match within 1 ULP.
        // ====================================================================
        $display("\nTest 7: Incremental interpolation accuracy");
        fb_width_log2  = 4'd9;
        fb_height_log2 = 4'd9;
        pixel_count = 0;

        // Triangle: V0=(10,10), V1=(30,10), V2=(20,30) -- small, fully on-screen
        v0_x = 16'd160;   // 10 << 4
        v0_y = 16'd160;   // 10 << 4
        v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;   // R=255, G=0, B=0, A=0
        v0_color1 = 32'h00000000;
        v0_uv0 = {16'h0000, 16'h0000};  // UV0=(0.0, 0.0)
        v0_uv1 = 32'h00000000;
        v0_q = 16'h1000;   // Q = 1.0 in Q3.12

        v1_x = 16'd480;   // 30 << 4
        v1_y = 16'd160;   // 10 << 4
        v1_z = 16'h3000;
        v1_color0 = 32'h00FF0000;   // R=0, G=255, B=0, A=0
        v1_color1 = 32'h00000000;
        v1_uv0 = {16'h1000, 16'h0000};  // UV0=(1.0, 0.0)
        v1_uv1 = 32'h00000000;
        v1_q = 16'h1000;

        v2_x = 16'd320;   // 20 << 4
        v2_y = 16'd480;   // 30 << 4
        v2_z = 16'h2000;
        v2_color0 = 32'h0000FF00;   // R=0, G=0, B=255, A=0
        v2_color1 = 32'h00000000;
        v2_uv0 = {16'h0000, 16'h1000};  // UV0=(0.0, 1.0)
        v2_uv1 = 32'h00000000;
        v2_q = 16'h2000;   // Q = 2.0 in Q3.12

        // 2*area = |(30-10)*(30-10)-(20-10)*(10-10)| = |20*20-10*0| = 400
        // inv_area = 65536/400 = 163.84 ~ 164 = 0x00A4
        inv_area = 16'h00A4;

        // Submit the triangle and collect fragments
        frag_ready = 1;
        submit_triangle_and_wait;
        $display("  Interpolation test completed, fragments=%0d", pixel_count);

        // After rasterization, compute reference values for the first fragment
        // position.  The rasterizer walks from bbox_min, so the first inside
        // pixel should be at or near vertex V0.  We verify that the DUT's
        // internal derivative registers match our reference computation.
        //
        // The rasterizer latches edge coefficients in SETUP state:
        //   edge1_A = y2 - y0 = 30 - 10 = 20
        //   edge1_B = x0 - x2 = 10 - 20 = -10
        //   edge2_A = y0 - y1 = 10 - 10 = 0
        //   edge2_B = x1 - x0 = 30 - 10 = 20
        //
        // Reference color0 R derivative dx:
        //   d10 = c0_r1 - c0_r0 = 0 - 255 = -255
        //   d20 = c0_r2 - c0_r0 = 0 - 255 = -255
        //   raw = (-255 * 20) + (-255 * 0) = -5100
        //   scl = -5100 * 164 = -836400
        //   dx  = -836400 >>> 16 = -12 (truncated)
        begin : interp_check
            reg signed [10:0] ref_e1A, ref_e1B, ref_e2A, ref_e2B;
            reg signed [31:0] ref_c0r_dx, ref_c0r_dy;
            reg signed [31:0] ref_c0g_dx, ref_c0g_dy;
            reg signed [31:0] ref_c0b_dx, ref_c0b_dy;
            reg signed [31:0] ref_z_dx, ref_z_dy;
            reg signed [31:0] ref_uv0u_dx, ref_uv0u_dy;
            reg signed [31:0] ref_uv0v_dx, ref_uv0v_dy;
            reg signed [31:0] ref_q_dx, ref_q_dy;
            integer interp_fail;

            // Edge coefficients from rasterizer (latched during SETUP)
            // Using pixel coordinates: x0=10, y0=10, x1=30, y1=10, x2=20, y2=30
            ref_e1A = $signed(11'd30) - $signed(11'd10);  // y2 - y0 = 20
            ref_e1B = $signed(11'd10) - $signed(11'd20);  // x0 - x2 = -10
            ref_e2A = $signed(11'd10) - $signed(11'd10);  // y0 - y1 = 0
            ref_e2B = $signed(11'd30) - $signed(11'd10);  // x1 - x0 = 20

            // Color0 R: f0=255, f1=0, f2=0
            ref_c0r_dx = ref_deriv_8bit(8'd255, 8'd0, 8'd0, ref_e1A, ref_e2A, 16'h00A4);
            ref_c0r_dy = ref_deriv_8bit(8'd255, 8'd0, 8'd0, ref_e1B, ref_e2B, 16'h00A4);

            // Color0 G: f0=0, f1=255, f2=0
            ref_c0g_dx = ref_deriv_8bit(8'd0, 8'd255, 8'd0, ref_e1A, ref_e2A, 16'h00A4);
            ref_c0g_dy = ref_deriv_8bit(8'd0, 8'd255, 8'd0, ref_e1B, ref_e2B, 16'h00A4);

            // Color0 B: f0=0, f1=0, f2=255
            ref_c0b_dx = ref_deriv_8bit(8'd0, 8'd0, 8'd255, ref_e1A, ref_e2A, 16'h00A4);
            ref_c0b_dy = ref_deriv_8bit(8'd0, 8'd0, 8'd255, ref_e1B, ref_e2B, 16'h00A4);

            // Z: z0=0x1000, z1=0x3000, z2=0x2000
            ref_z_dx = ref_deriv_16bit(
                $signed({1'b0, 16'h3000}) - $signed({1'b0, 16'h1000}),
                $signed({1'b0, 16'h2000}) - $signed({1'b0, 16'h1000}),
                ref_e1A, ref_e2A, 16'h00A4);
            ref_z_dy = ref_deriv_16bit(
                $signed({1'b0, 16'h3000}) - $signed({1'b0, 16'h1000}),
                $signed({1'b0, 16'h2000}) - $signed({1'b0, 16'h1000}),
                ref_e1B, ref_e2B, 16'h00A4);

            // UV reference values are Q4.12 (16-bit signed: sign [15], integer [14:12], fractional [11:0])
            // per UNIT-005 fragment bus spec and fp_types_pkg.sv q4_12_t typedef.

            // UV0 U: u0=0x0000, u1=0x1000, u2=0x0000
            ref_uv0u_dx = ref_deriv_16bit(
                {1'b0, 16'h1000} - {1'b0, 16'h0000},
                {1'b0, 16'h0000} - {1'b0, 16'h0000},
                ref_e1A, ref_e2A, 16'h00A4);
            ref_uv0u_dy = ref_deriv_16bit(
                {1'b0, 16'h1000} - {1'b0, 16'h0000},
                {1'b0, 16'h0000} - {1'b0, 16'h0000},
                ref_e1B, ref_e2B, 16'h00A4);

            // UV0 V: v0=0x0000, v1=0x0000, v2=0x1000
            ref_uv0v_dx = ref_deriv_16bit(
                {1'b0, 16'h0000} - {1'b0, 16'h0000},
                {1'b0, 16'h1000} - {1'b0, 16'h0000},
                ref_e1A, ref_e2A, 16'h00A4);
            ref_uv0v_dy = ref_deriv_16bit(
                {1'b0, 16'h0000} - {1'b0, 16'h0000},
                {1'b0, 16'h1000} - {1'b0, 16'h0000},
                ref_e1B, ref_e2B, 16'h00A4);

            // Q: q0=0x1000, q1=0x1000, q2=0x2000
            ref_q_dx = ref_deriv_16bit(
                $signed({1'b0, 16'h1000}) - $signed({1'b0, 16'h1000}),
                $signed({1'b0, 16'h2000}) - $signed({1'b0, 16'h1000}),
                ref_e1A, ref_e2A, 16'h00A4);
            ref_q_dy = ref_deriv_16bit(
                $signed({1'b0, 16'h1000}) - $signed({1'b0, 16'h1000}),
                $signed({1'b0, 16'h2000}) - $signed({1'b0, 16'h1000}),
                ref_e1B, ref_e2B, 16'h00A4);

            interp_fail = 0;

            $display("  Derivative verification (DUT vs reference):");

            // Check color0 R dx
            $display("    c0r_dx: DUT=%0d, ref=%0d", dut.c0r_dx, ref_c0r_dx);
            if (dut.c0r_dx == ref_c0r_dx) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: c0r_dx mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check color0 R dy
            $display("    c0r_dy: DUT=%0d, ref=%0d", dut.c0r_dy, ref_c0r_dy);
            if (dut.c0r_dy == ref_c0r_dy) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: c0r_dy mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check color0 G dx
            $display("    c0g_dx: DUT=%0d, ref=%0d", dut.c0g_dx, ref_c0g_dx);
            if (dut.c0g_dx == ref_c0g_dx) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: c0g_dx mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check color0 G dy
            $display("    c0g_dy: DUT=%0d, ref=%0d", dut.c0g_dy, ref_c0g_dy);
            if (dut.c0g_dy == ref_c0g_dy) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: c0g_dy mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check color0 B dx
            $display("    c0b_dx: DUT=%0d, ref=%0d", dut.c0b_dx, ref_c0b_dx);
            if (dut.c0b_dx == ref_c0b_dx) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: c0b_dx mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check color0 B dy
            $display("    c0b_dy: DUT=%0d, ref=%0d", dut.c0b_dy, ref_c0b_dy);
            if (dut.c0b_dy == ref_c0b_dy) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: c0b_dy mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check Z dx
            $display("    z_dx:   DUT=%0d, ref=%0d", dut.z_dx, ref_z_dx);
            if (dut.z_dx == ref_z_dx) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: z_dx mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check Z dy
            $display("    z_dy:   DUT=%0d, ref=%0d", dut.z_dy, ref_z_dy);
            if (dut.z_dy == ref_z_dy) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: z_dy mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check UV0 U dx (Q4.12)
            $display("    uv0u_dx (Q4.12): DUT=%0d, ref=%0d", dut.uv0u_dx, ref_uv0u_dx);
            if (dut.uv0u_dx == ref_uv0u_dx) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: uv0u_dx (Q4.12) mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check UV0 U dy (Q4.12)
            $display("    uv0u_dy (Q4.12): DUT=%0d, ref=%0d", dut.uv0u_dy, ref_uv0u_dy);
            if (dut.uv0u_dy == ref_uv0u_dy) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: uv0u_dy (Q4.12) mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check UV0 V dx (Q4.12)
            $display("    uv0v_dx (Q4.12): DUT=%0d, ref=%0d", dut.uv0v_dx, ref_uv0v_dx);
            if (dut.uv0v_dx == ref_uv0v_dx) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: uv0v_dx (Q4.12) mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check UV0 V dy (Q4.12)
            $display("    uv0v_dy (Q4.12): DUT=%0d, ref=%0d", dut.uv0v_dy, ref_uv0v_dy);
            if (dut.uv0v_dy == ref_uv0v_dy) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: uv0v_dy (Q4.12) mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check Q dx
            $display("    q_dx:   DUT=%0d, ref=%0d", dut.q_dx, ref_q_dx);
            if (dut.q_dx == ref_q_dx) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: q_dx mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            // Check Q dy
            $display("    q_dy:   DUT=%0d, ref=%0d", dut.q_dy, ref_q_dy);
            if (dut.q_dy == ref_q_dy) begin
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("    FAIL: q_dy mismatch");
                test_fail_count = test_fail_count + 1;
                interp_fail = 1;
            end

            if (interp_fail == 0) begin
                $display("  PASS: All derivative registers match reference model (UV0, UV1 (Q4.12))");
            end else begin
                $display("  FAIL: One or more derivative registers differ from reference (UV0, UV1 (Q4.12))");
            end
        end

        repeat(20) @(posedge clk);

        // ====================================================================
        // Test 8: Winding order (VER-001 step 7)
        // Submit the same triangle in CCW and CW winding order.
        // Verify that edge function signs are consistent with the expected
        // winding convention and that fragment emission occurs for the
        // correct winding.
        // ====================================================================
        $display("\nTest 8: Winding order test");
        fb_width_log2  = 4'd9;
        fb_height_log2 = 4'd9;

        // --- 8a: Counter-clockwise winding (V0-V1-V2 forms CCW) ---
        $display("  8a: Counter-clockwise winding");
        pixel_count = 0;

        // V0=(10,10), V1=(30,10), V2=(20,30) -- CCW when Y increases downward
        v0_x = 16'd160;  v0_y = 16'd160;  v0_z = 16'h1000;
        v0_color0 = 32'hFF000000;
        set_default_attrs;

        v1_x = 16'd480;  v1_y = 16'd160;  v1_z = 16'h2000;
        v1_color0 = 32'h00FF0000;

        v2_x = 16'd320;  v2_y = 16'd480;  v2_z = 16'h3000;
        v2_color0 = 32'h0000FF00;

        inv_area = 16'h00A4;

        submit_triangle_and_wait;
        $display("    CCW fragments=%0d", pixel_count);

        begin : winding_ccw
            integer ccw_count;
            ccw_count = pixel_count;

            // --- 8b: Clockwise winding (swap V1 and V2) ---
            $display("  8b: Clockwise winding (V1 and V2 swapped)");
            pixel_count = 0;

            // V0=(10,10), V1=(20,30), V2=(30,10) -- CW
            v0_x = 16'd160;  v0_y = 16'd160;  v0_z = 16'h1000;
            v0_color0 = 32'hFF000000;
            set_default_attrs;

            v1_x = 16'd320;  v1_y = 16'd480;  v1_z = 16'h3000;
            v1_color0 = 32'h0000FF00;

            v2_x = 16'd480;  v2_y = 16'd160;  v2_z = 16'h2000;
            v2_color0 = 32'h00FF0000;

            inv_area = 16'h00A4;

            submit_triangle_and_wait;
            $display("    CW fragments=%0d", pixel_count);

            // The edge function convention should produce fragments for one
            // winding and not the other (or produce the same count for both
            // if the rasterizer is winding-agnostic with abs(area)).
            // At minimum, verify that both triangle submissions complete
            // successfully and that the fragment counts are consistent.
            if (ccw_count > 0 || pixel_count > 0) begin
                $display("  PASS: Winding order test -- CCW=%0d, CW=%0d fragments", ccw_count, pixel_count);
                test_pass_count = test_pass_count + 1;
            end else begin
                $display("  FAIL: Neither winding order produced fragments");
                test_fail_count = test_fail_count + 1;
            end

            // Edge function signs should be inverted between CW and CCW.
            // Check that edge0_A differs in sign (or both are zero for
            // horizontal edges).
            $display("    Edge0_A (after CW): %0d", dut.edge0_A);
        end

        repeat(20) @(posedge clk);

        // ====================================================================
        // Summary
        // ====================================================================
        $display("\n=== Rasterizer Test Summary ===");
        $display("  Passed: %0d", test_pass_count);
        $display("  Failed: %0d", test_fail_count);
        $display("  Total fragments emitted: %0d", total_frag_count);

        if (test_fail_count == 0) begin
            $display("RESULT: PASS");
        end else begin
            $display("RESULT: FAIL");
        end

        $display("=== Rasterizer Test Completed ===");
        $finish;
    end

    // Timeout watchdog
    initial begin
        #20000000;  // 20ms timeout (increased for interpolation and winding tests)
        $display("\nERROR: Timeout - simulation ran too long");
        $finish;
    end

endmodule
